
module test_Huang();
    initial begin
        $display("Hello, Huang");
        end
endmodule