
module Hello_World;

initial begin
    $display("Hello, World");
end

endmodule