module led_test(input key_in,output led_out);
assign led_out=~key_in;

endmodule